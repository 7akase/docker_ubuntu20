class  extends ;
`uvm_component_utils()

function new(string name, uvm_component parent);
    super.new(name, parent);
endfunction

endclass