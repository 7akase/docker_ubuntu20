`define CBLK    $write("%c[1;30m",27);
`define CRED    $write("%c[1;31m",27);
`define CGREEN  $write("%c[1;32m",27);
`define CBLUE   $write("%c[1;34m",27);
`define CEND    $write("%c[0m",27);