class  extends ;
`uvm_object_utils()

function new(string name="");
    super.new(name);
endfunction

endclass