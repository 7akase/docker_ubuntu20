class aaa extends uvm_object;
    `uvm_object_utils()

    function new(string name="");
        super.new(name);
    endfunction

    // extern task pre_body();
    // extern task body();
    // extern task post_body();
endclass
